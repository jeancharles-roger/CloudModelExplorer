
cdl test1 is {
	main is {event {send "hello" to {process}1}}
}
