
cdl test1 is {
	main is {
		event {send "hello" to {process}1} ||
		event {send "hello" to {process}2} ||
		event {send "hello" to {process}3} ||
		event {send "hello" to {process}4}
	}
}
